`timescale 1ns / 1ps
////////////////////////////////////////////////////////
// Assignment 6 - CS31001
// Implementing Diff Operation
// Team Details - 
// Kushaz Sehgal - 20CS30030
// Jay Kumar Thakur - 20CS30024
////////////////////////////////////////////////////////

module Diff(
    input [31:0] a,
    input [31:0] b,
    output [31:0] c
);

    wire [31:0] xor_ab, index_num,carry_buffer; 
    assign xor_ab = a^b;

    Adder_32_bit minus_1(.a(xor_ab),.b(32'b11111111111111111111111111111111),.c_in(32'b00000000000000000000000000000000),.sum(index_num),.c_out(carry_buffer))
    
    always @(*) begin
        case (index_num)
            32'b00000000000000000000000000000001 : c = 32'd1 
            32'b00000000000000000000000000000010 : c = 32'd1 
            32'b00000000000000000000000000000100 : c = 32'd1 
            32'b00000000000000000000000000001000 : c = 32'd1 
            32'b00000000000000000000000000010000 : c = 32'd1 
            32'b00000000000000000000000000100000 : c = 32'd1 
            32'b00000000000000000000000001000000 : c = 32'd1 
            32'b00000000000000000000000010000000 : c = 32'd1
            32'b00000000000000000000000100000000 : c = 32'd1 
            32'b00000000000000000000001000000000 : c = 32'd1 
            32'b00000000000000000000010000000000 : c = 32'd1 
            32'b00000000000000000000100000000000 : c = 32'd1 
            32'b00000000000000000001000000000000 : c = 32'd1 
            32'b00000000000000000010000000000000 : c = 32'd1 
            32'b00000000000000000100000000000000 : c = 32'd1 
            32'b00000000000000001000000000000000 : c = 32'd1
            32'b00000000000000010000000000000000 : c = 32'd1 
            32'b00000000000000100000000000000000 : c = 32'd1 
            32'b00000000000001000000000000000000 : c = 32'd1 
            32'b00000000000010000000000000000000 : c = 32'd1 
            32'b00000000000100000000000000000000 : c = 32'd1 
            32'b00000000001000000000000000000000 : c = 32'd1 
            32'b00000000010000000000000000000000 : c = 32'd1 
            32'b00000000100000000000000000000000 : c = 32'd1
            32'b00000001000000000000000000000000 : c = 32'd1 
            32'b00000010000000000000000000000000 : c = 32'd1 
            32'b00000100000000000000000000000000 : c = 32'd1 
            32'b00001000000000000000000000000000 : c = 32'd1 
            32'b00010000000000000000000000000000 : c = 32'd1 
            32'b00100000000000000000000000000000 : c = 32'd1 
            32'b01000000000000000000000000000000 : c = 32'd1 
            32'b10000000000000000000000000000000 : c = 32'd1 
            default : c = 32'd0
    end
endmodule
