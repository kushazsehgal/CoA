module not(o, i):
    input i;
    ouput o;
    not(o, i);
endmodule